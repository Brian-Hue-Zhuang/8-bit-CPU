module machine (
    input logic clk, rst
);
    logic [7:0] data_bus;
    tri [7:0] bus;
    logic wEN, wEN, clk;
endmodule